.title KiCad schematic
.include "C:/AE/LP38693/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/LP38693/_models/LP38693_ADJ_TRANS.lib"
.include "C:/AE/LP38693/_models/PCF1C101MCL1GS_v100.lib"
.include "C:/AE/LP38693/_models/PCF1E100MCL1GS_v100.lib"
XU4 /VOUT 0 PCF1C101MCL1GS
R2 /VOUT /VADJ {RADJ}
R3 /VADJ 0 {RREF}
XU3 /VIN /VADJ /EN /VOUT 0 LP38693_ADJ_TRANS
XU5 /VOUT 0 C2012X7R2A104K125AA_p
I1 /VOUT 0 {ILOAD}
R1 /VIN /EN {REN}
V1 /VIN 0 {VSOURCE}
XU1 /VIN 0 PCF1E100MCL1GS
XU2 /VIN 0 C2012X7R2A104K125AA_p
.end
